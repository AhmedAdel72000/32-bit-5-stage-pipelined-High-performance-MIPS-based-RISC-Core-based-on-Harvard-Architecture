module ADD (INPUT1 , INPUT2 , ADDRESULT);
input [31:0] INPUT1 , INPUT2 ;
output ADDRESULT ;
assign ADDRESULT = INPUT1 + INPUT2 ;
endmodule
